library verilog;
use verilog.vl_types.all;
entity clock_vlg_check_tst is
    port(
        clk             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end clock_vlg_check_tst;
