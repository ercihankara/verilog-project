library verilog;
use verilog.vl_types.all;
entity son_vlg_vec_tst is
end son_vlg_vec_tst;
