library verilog;
use verilog.vl_types.all;
entity take_in_in_vlg_vec_tst is
end take_in_in_vlg_vec_tst;
