library verilog;
use verilog.vl_types.all;
entity read_new_vlg_vec_tst is
end read_new_vlg_vec_tst;
