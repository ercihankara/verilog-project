library verilog;
use verilog.vl_types.all;
entity read_vlg_vec_tst is
end read_vlg_vec_tst;
